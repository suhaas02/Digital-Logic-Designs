module priority_dec
